Iniciando teste da Control Unit...
=================================
Tempo                   10: Opcode=000000 (R-type) | RegDst=1, Branch=0, MemRead=0, MemtoReg=0, ALUOp=10, MemWrite=0, ALUSrc=0, RegWrite=1
Tempo                   20: Opcode=100011 (lw)     | RegDst=0, Branch=0, MemRead=1, MemtoReg=1, ALUOp=00, MemWrite=0, ALUSrc=1, RegWrite=1
Tempo                   30: Opcode=101011 (sw)     | RegDst=0, Branch=0, MemRead=0, MemtoReg=1, ALUOp=00, MemWrite=1, ALUSrc=1, RegWrite=0
Tempo                   40: Opcode=000100 (beq)    | RegDst=0, Branch=1, MemRead=0, MemtoReg=1, ALUOp=01, MemWrite=0, ALUSrc=0, RegWrite=0
Tempo                   50: Opcode=001000 (addi)   | RegDst=0, Branch=0, MemRead=0, MemtoReg=0, ALUOp=00, MemWrite=0, ALUSrc=1, RegWrite=1
Tempo                   60: Opcode=111111 (inválido)| RegDst=0, Branch=0, MemRead=0, MemtoReg=0, ALUOp=00, MemWrite=0, ALUSrc=0, RegWrite=0
=================================
Teste da Control Unit concluído com sucesso!
