
Tempo                    0: opcode=000000 | RegDst=1, Branch=0, MemRead=0, MemtoReg=0, ALUOp=10, MemWrite=0, ALUSrc=0, RegWrite=1
Tempo                   30: opcode=100011 | RegDst=0, Branch=0, MemRead=1, MemtoReg=1, ALUOp=00, MemWrite=0, ALUSrc=1, RegWrite=1
Tempo                   50: opcode=101011 | RegDst=0, Branch=0, MemRead=0, MemtoReg=1, ALUOp=00, MemWrite=1, ALUSrc=1, RegWrite=0
Tempo                   70: opcode=000100 | RegDst=0, Branch=1, MemRead=0, MemtoReg=1, ALUOp=01, MemWrite=0, ALUSrc=0, RegWrite=0
Tempo                   90: opcode=001000 | RegDst=0, Branch=0, MemRead=0, MemtoReg=0, ALUOp=00, MemWrite=0, ALUSrc=1, RegWrite=1
Tempo                  110: opcode=111111 | RegDst=0, Branch=0, MemRead=0, MemtoReg=0, ALUOp=00, MemWrite=0, ALUSrc=0, RegWrite=0
Testes concluídos!
