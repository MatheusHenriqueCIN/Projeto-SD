Iniciando teste da DataMemory...
=================================
[MEM WRITE] Addr: 00000004 : Data: abcd1234
[MEM READ] Addr: 00000004 : Data: abcd1234
[MEM WRITE] Addr: 00000ffc : Data: ffffffff
[MEM READ] Addr: 00000ffc : Data: ffffffff
[MEM READ ERROR] Endereço 00001000 fora dos limites!
=================================
Teste da DataMemory concluído!
