Iniciando teste do PC Branch...
=================================

Teste 1 - PC+4: 0x00001004, Imm: 0x00000001 -> PCBranch: 0x00001008 (Esperado: 0x00001008)
Teste 2 - PC+4: 0x00002008, Imm: 0x00000100 -> PCBranch: 0x00002408 (Esperado: 0x00002408)
Teste 3 - PC+4: 0x0000300c, Imm: 0xfffffffc -> PCBranch: 0x00002ffc (Esperado: 0x00002ffc)
Teste 4 - PC+4: 0x00004010, Imm: 0x00000000 -> PCBranch: 0x00004010 (Esperado: 0x00004010)
Teste 5 - PC+4: 0x7ffffffc, Imm: 0x3fffffff -> PCBranch: 0x7ffffff8 (Esperado: 0x7ffffff8)

=================================
Teste do PC Branch concluído com sucesso!
